package aes_const;
  timeunit 1ns;
  timeprecision 1ps;

  // parameter Nb = 4;
  // parameter Nk = 4;
  // parameter Nr = 10;
  //
  // parameter [127:0] key = 128'h2b7e151628aed2a6abf7158809cf4f3c;
  // parameter [127:0] data = 128'h0;

  // parameter Nb = 4;
  // parameter Nk = 6;
  // parameter Nr = 12;
  //
  // parameter [191:0] key = 192'h8e73b0f7da0e6452c810f32b809079e562f8ead2522c6b7b;
  // parameter [127:0] data = 128'h0;

  // parameter Nb = 4;
  // parameter Nk = 8;
  // parameter Nr = 14;
  //
  // parameter [255:0] key = 256'h603deb1015ca71be2b73aef0857d77811f352c073b6108d72d9810a30914dff4;
  // parameter [127:0] data = 128'h0;

  parameter Nb = 4;
  parameter Nk = 4;
  parameter Nr = 10;

  parameter [127:0] key = 128'h2b7e151628aed2a6abf7158809cf4f3c;
  parameter [127:0] data = 128'h03243f6a8885a308d313198a2e0370734;

endpackage
