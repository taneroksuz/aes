package aes_const;
	timeunit 1ns;
	timeprecision 1ps;

  localparam  Nb = 4;
  localparam  Nk = 4;
  localparam  Nr = 10;

endpackage
